`define DELAY 20
module _32bit_adder_testbench();
reg [31:0] a, b;

wire [31:0] s;


_32bit_adder a1(s,a,b);

initial begin

a = 32'b10000000000000000000000000000000; b = 32'b10000000000000000000000000000000;
#`DELAY;
a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000001;
#`DELAY;
a = 32'b01000000000000000000000000000000; b = 32'b01000000000000000000000000000001;
#`DELAY;
a = 32'b00000000000000000000000000010000; b = 32'b00000000000000000000000000001001;
end
 
 
initial
begin
$monitor("time = %2d, out=%32b", $time, s);
end
 
endmodule