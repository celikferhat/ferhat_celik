`define DELAY 20
module _32bit_alu_testbench(); 
reg [31:0]a, b;
reg [2:0]select;
wire [31:0] out;
wire v , z , carry_out;
alu32 al(out,v,z,carry_out, a, b, select);

initial begin

// AND
a = 32'b00100100001010001110000000000100; b = 32'b00100100001010001110000000011110; select = 3'b000;
#`DELAY;
a = 32'b11111111111111111111111111111111; b = 32'b00000000000000000000000000000001; select = 3'b000;
#`DELAY;
a = 32'b10111010111101010111111110111100; b = 32'b10101111100101011111110101011110; select = 3'b000;
#`DELAY;
// OR
a = 32'b01000000000000000000000000000001; b = 32'b11000000000000000000000000000100; select = 3'b001;
#`DELAY;
a = 32'b11111111111111111111111111111111; b = 32'b00000000000000000000000000000001; select = 3'b001;
#`DELAY;
a = 32'b01000010000000001010110100000001; b = 32'b11010010111101111101010000000100; select = 3'b001;
#`DELAY;
// ADD
a = 32'b01100011111111011010100000011100; b = 32'b10000010000010111000000000011000; select = 3'b010;
#`DELAY;
a = 32'b01000000000111010110000000000001; b = 32'b01111100000000000000011100000100; select = 3'b010;
#`DELAY;
a = 32'b11000000000000000000000000000001; b = 32'b01000000000000000000000000000100; select = 3'b010;
#`DELAY;

// SUBSTRACT
a = 32'b00000000000000000000000000000001; b = 32'b00000000000000000000000000000010; select = 3'b110;
#`DELAY;
a = 32'b01110110100000000000000000000001; b = 32'b00011011011111010111000000000100; select = 3'b110;
#`DELAY;
a = 32'b11000000000000000000000000000001; b = 32'b10000001111011011000000000000100; select = 3'b110;
#`DELAY;

// SLT
a = 32'b01110101010101111111010101010101; b = 32'b11010111110110101111101010101010; select = 3'b111;
#`DELAY;
a = 32'b11000000000000000000000000000001; b = 32'b11000000000000000000000000000100; select = 3'b111;
#`DELAY;
a = 32'b01110101111101011111110000000001; b = 32'b10011101111101110000000000000100; select = 3'b111;
#`DELAY;
a = 32'b01110101111101011111110000000001; b = 32'b10011101111101110000000000000100; select = 3'b011;
#`DELAY;
end
 
 
initial
begin
$monitor("time = %2d, Input1 = %32b, Input2 = %32b, select=%3b, out=%32b ,v=%1b ,z=%1b, carry_out=%1b", $time, a, b, select, out,v,z,carry_out);
end
 
endmodule